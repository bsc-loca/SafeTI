-----------------------------------------------------------------------------   
-- Entity:      axi4_manager
-- File:        axi4_manager.vhd
-- Author:      Francisco Javier Fuentes Diaz (BSC-CNS)
-- Description: AXI4 FULL Manager entity.
------------------------------------------------------------------------------ 
--  Changelog:
--              - v0.8.9  WIP.
--                The interface has been reworked, in such a way where the logic has been split 
--                between handshake (hs) and burst (burst) state machines, in order to allow granting 
--                transactions on the BM side even when a transaction are ongoing at the AXI side.
--                This means that the interface may now generate requests at the AXI side during a 
--                burst transfer of the previous BM transaction.
--                If the burst is granted, that burst will not initiate until the ongoing one ends.
--                Enabling "injector_mode" allows to simulate the BM signaling without really making 
--                any data transfer between the BM component and the interface. Read data is discarded 
--                and write data is zeroed.
--                Due to some bugs that have been detected, this version is WIP. 
--
--              - v0.8.6  May  5, 2022.
--                Added input signals for setting the AXI burst parameters as fixed address 
--                transactions, CACHE and PROT, so they can be configured by the BM component.
--                The Injector_implementation option has been dropped, since the functionality 
--                did not save particulary many resources while not being that useful if the BM 
--                component scales correctly with dbits.
--
--              - v0.8.5  Mar 29, 2022.
--                Now the rd.bm_valid is asserted correctly on discarded data read transactions
--                due to Injector_implementation being TRUE.
--                All AXI parametrizable variables, as bus widths, have been moved to generics.
--                This, while making easier the integration of the interface, it also has 
--                expanded the bus widths to the maximum allowed by the protocol, in order to 
--                accomodate such cases. However, the synthesis tool should remove unnused wiring.
--
--              - v0.8.2  Mar 11, 2022.
--                Configurable parameters of the number of FIFO registers and injector 
--                mode have been moved as generics, allowing multiple instances with 
--                different properties. AXI infrastructure properties are still general, thou.
--
--              - v0.8.1  Mar  1, 2022.
--                I/O types for the BM component have been renamed to bm_miso and
--                bm_mosi, while the AXI I/O types have been renamed axi4_miso and
--                axi4_mosi. In this aspect, the design perspective is that the BM
--                component is the "Manager" for the interface, while the interface is 
--                the subordinate for the BM component. Thus, the BM componente outputs 
--                MOSI signals to the interface, and the interface outputs MISO signals 
--                to the BM component.
--                Bug solved where the write strobe would be incorrect at the last beat of  
--                the burst if the beat was not transmited (w_ready = 1) on that cycle.
--                Modifications have been made to achieve synthesis in isolated module mode.
--
--              - v0.8    Feb 25, 2022. 
--                First deliver of the AXI Manager interface as a working module.
--                It has passed manual debugging. There may be errors not found, 
--                specially on write transactions. Contact the author through GitLab 
--                opening an issue ticket specifying the request data and the problem.
--                Synthesis optimization is yet to be done.
--
------------------------------------------------------------------------------ 

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library safety;
use safety.axi4_pkg.all; -- <- It contains the configuration of the interface.

-----------------------------------------------------------------------------
-- AXI4 FULL Manager - bus manager bridge
--
-- Manager interface features:
--
-- - Only INC burst mode is available and every burst generated use all AXI data lanes available per beat.
-- - Full support for unaligned address requests. This includes even if two subordinates are accessed in a 
--   single transaction request.
-- - Number of bytes per BM transaction requests allowed is 4096 (encoded as 0xFFF).
-- - BM done output flag assertion at the end of every transaction on its appropiated bus (reads or writes).
-- - Extensible BM component and AXI data buses width 8, 16, 32, 64, 128, 256, 512 and 1024 bits (read 
--   further considerations on integration of the interface for limitations).
-- - Continuous data transmission if there's enough data supply throughput from the least data bus bottleneck.
--
--
-- Manager interface and considerations during integration:
--
-- - DATA_WIDTH >= dbits. The AXI data bus width must be greater or equal to the BM data bus.
--
-- - BM size requests <= 4096 (4kB, limited by AXI4 addressing rule). The maximum number of bytes 
--   per BM transaction is 4096 (encoded as 0xFFF).
--
-- - Little endian data structure. Higher bit position links to higher memory positions.
--
-- - Only INC burst mode is implemented. This is the mode where the addressing increases every beat 
--   at AXI data width bytes steps on the AXI side.
--
-- - Unaligned access by BM requests are supported through aligning the address with AXI data bus width,
--   while delivering only the requested data on read transactions and using the write strobe on AXI 
--   write transactions.
--
-- - The Manager only execute bursts with the AXI size that use the whole AXI data bus width.
--
-- - This interface requires the signaling of the last AXI beat to be at the correct beat on read 
--   transactions, or unrequested data could be read instead of the requested.
--
-- - The interface may send control and data when the valid flag is not asserted. These signals 
--   must be discarded since the valid flag is low.
--
--
-- This AXI4 Manager interface translates and manage the requests made by the BM component,
-- using the BM input and output buses, to the AXI4 network, using the AXI4 input and output buses.
--
-- The BM component has an opaque vision of what the interface requests to the AXI network, since 
-- it only receives the data that it has been requested. Be it requests with unaligned or even to multiple 
-- subordinates access (only 2 as maximum), the interface filters it to deliver only the requested data.
-- 
-- Most I/O ports are buffered on registers to promote higher maximum frequency of operation at 
-- implementation, with minimum logic between register and BM or AXI bus. In any case, there is not
-- a direct I/O path that could greatly impact the fMAX once the interface is integrated on the project.
-- 
-- If the BM request implies access to two different subordinates, the Manager interface will generate two 
-- batches of data that are distribuited in one or multiple bursts each, with the appropiated addressing 
-- and burst length (number of beats in the burst) for each burst). Multiple bursts for the same batch
-- depends on the AXI data bus width, since implemenations with an AXI data bus width lower than 128 bits 
-- require multiple bursts to the same subordinate to be able to access the 4kB of data (4096 addresses) 
-- it can allocate (limit listed by the AXI4 protocol).
-- 
-- 
-----------------------------------------------------------------------------

entity axi4_manager is
  generic (
    -- AXI Manager configuration
    ID_R_WIDTH      : integer range  0 to   32  := 4;       -- AXI ID's bus width.
    ID_W_WIDTH      : integer range  0 to   32  := 4;       -- AXI ID's bus width.
    ADDR_WIDTH      : integer range 12 to   64  := 32;      -- AXI address bus width. (Tested only for 32 bits)
    DATA_WIDTH      : integer range  8 to 1024  := 128;     -- AXI data bus width. [Only power of 2s are allowed]
    axi_id          : integer range  0 to 32**2-1 := 0;     -- AXI manager burst index [Must be < ID_X_WIDTH**2-1]
    injector_mode   : boolean                   := TRUE;   -- Simulate read BM transfers to save on footprint

    -- Bus Manager (BM) configuration
    dbits           : integer range  8 to 1024  := 32;      -- BM data bus width [Only power of 2s are allowed and <= AXI_DATA_WIDTH]

    -- Interface configuration
    rd_n_fifo_regs  : integer range  2 to  256  := 2;       -- Number of FIFO registers to use at AXI read transactions.  [Only power of 2s are allowed]
    wr_n_fifo_regs  : integer range  2 to  256  := 2;       -- Number of FIFO registers to use at AXI write transactions. [Only power of 2s are allowed]
    ASYNC_RST       : boolean                   := FALSE    -- Allow asynchronous reset
  );
  port (
    rstn                      : in  std_ulogic; -- Reset
    clk                       : in  std_ulogic; -- Clock
    -- AXI interface signals
    axi4mi                    : in  axi4_miso;  -- AXI4 manager input 
    axi4mo                    : out axi4_mosi;  -- AXI4 manager output
    -- BM component signals
    bm_in                     : in  bm_mosi;    -- BM interface input
    bm_out                    : out bm_miso     -- BM interface output
  );
end entity axi4_manager;

architecture rtl of axi4_manager is
  -----------------------------------------------------------------------------
  -- Constant declaration
  -----------------------------------------------------------------------------

    -- Parametric constants
    constant DBITS_DATA_BYTE  : integer := log_2(dbits/8);      -- Number of bits required to address the BM data bus bytes.
    constant AXI4_DATA_BYTE   : integer := log_2(DATA_WIDTH/8); -- Number of bits required to address the AXI data bus bytes.
    constant MAX_BURST_BYTE   : integer := log_2(4096);         -- Number of bits required to address the maximum transfer size by the protocol.

    -- The Mult_bursts_subor flag indicates when TRUE that the implementation allows for the possible requirement of multiple bursts to the same 
    -- subordinate (same 4kB memory space) to satisfy the size requested by the BM component (maximum 4096 bytes, encoded as 0xFFF in bm_in.bm_size).
    constant Mult_bursts_subor: boolean := DATA_WIDTH < 128;

  -----------------------------------------------------------------------------
  -- Records and types
  -----------------------------------------------------------------------------
  --
  -- This interface, when idle, accepts read and write transaction requests from the BM bus, listening the starting address and the total 
  -- transfer size of the operation. This last must be lower or equal to 4096 and it is encoded as an unsigned integer decremented by one 
  -- respect the real size. So a bm_in.rd_data 0x000 means 1 byte transfer, and the maximum is 0xFFF that is 4096 bytes to transfer.
  --
  -- Once the request has been granted (deassert granting new requests for that type of transaction until finished), the interface processes 
  -- the control data to check if the total transfer surpasses the 4kB address boundary, splitting the transaction in two batches 
  -- in such situations. This is done to arrange the transfer sizes of the batches for the first and second AXI subordinates, having 
  -- each different 4kB address allocation spaces.
  -- 
  -- Then, the interface sets an AXI size mode to use the whole data bus width of the AXI side (DATA_WIDTH), computes the number of beats 
  -- (burst length) to satisfy the request transfer and aligns the address requested (bm_addr) with the AXI data bus width (DATA_WIDTH).
  -- In case a single burst is not enough to satisfy the transfer size for the subordinate in question, the maximum length will be set (256 beats).
  -- However, this can only happen at implementations that have an DATA_WIDTH < 128 bits. Thus, this is managed with the "Mult_bursts_subor"
  -- flag to only proceed with the correspondent checks to generate multiple bursts to the same subordinate in the implementation if it's the case.
  --
  -- Since the BM component may request access to an unaligned address respect the DATA_WIDTH slot, the interface rearrenges the data to only 
  -- transfer to the BM component the data from the address requested on read transactions and to start writting from the address requested using 
  -- the byte strobe (wr.axi_strobe) on write transactions, even though the AXI Manager interface may request access to more data bytes.
  --
  -- The interface depends on the assertion of the AXI last signal on the last beat of the burst on read transactions in order to stop the transfer. 
  -- Otherwise, the interface may read data from the AXI data bus that should not and may transfered to the BM component instead of the requested data.
  -- 
  --
  -- The following table summarizes the actions done at each stage of the operation in both and on each type of transaction:
  -- 
  -- IDLE     -> Accept new requests from BM component.
  -- CHECK_4kB-> Compute if 4KB address space overflow occurs calculating the ending address of the BM request.
  --             In the case it does, assert burst_4kb flag so a second data batch is processed after completing the first.
  --             Also, split the total byte size of the transfer in both first and last batches taking into account the 4kB boundary.
  --          RD:Register the number of bytes to transfer at the last BM transfer of the whole transaction. This value is used to generate
  --             the mask applied on this last BM transfer, so unrequested data is not sent to the BM component.
  -- PREPARE_HS->Set the AXI size mode to use the whole AXI data bus width (encoded as log2(DATA_WIDTH/8)). 
  --             Also, generate an aligned address with the DATA_WIDTH slot to be used at the AXI network handshake.
  --             Set the burst mode (at the moment, this interface does only apply INC bursts).
  --             Decide burst length (number of beats) taking into the number of bytes to transfer and the address requested.
  --             Assert the AX valid signal (X is R for read or W for write transactions) to process the handshake of the burst.
  -- HANDSHAKE-> Waits for a AXI X ready input signal assertion so the handshake is executed and the AXI transfer can start.
  -- TRANSFER -> On the end of a burst on both transaction types (read transactions require the assertion of the last beat input signal 
  --             by part of the subordinate on the correct beat), the interface will check if any more data must be requested to the 
  --             actual subordinate. In affirmative case, another burst will be generated with the leftover number of bytes to transfer
  --             and the appropiated address. However, if it's not the case, be it because the BM size request is low enough or the 
  --             AXI data bus width is greater than 64 bits (4kB access is achievable in a single burst), the interface will generate 
  --             another burst to the next subordinate (next 4kB address space) with the leftover size requested. On both cases, this means 
  --             to return to the PREPARE_HS state with a different bm_size and bm_addr. 
  --             Once there's not leftover data to be transfered, it returns to the idle state, accepting new requests.
  --          RD:Reads the AXI data bus and register it onto rd_burst.axi_data_buffer if the AXI network reports valid data.
  --             After each beat (AXI data bus read), a FIFO register loads the data buffer, while also setting the rd_burst.fifo_full flag 
  --             for that particular register and increments the FIFO index, so the next FIFO register loads another beat from the buffer.
  --             In the case where all FIFO registers are full, the interface stops the read on the AXI data bus by deasserting rd_burst.axi_ready.
  --          WR:Set the strobe bits for WRITE transaction in accordance with the bytes that must be written on this beat.
  --             Load into wr.axi_data_buffer the data stored on the FIFO register, while asserting the wr.axi_valid_data so a beat is 
  --             transfered to the AXI network on the next clock cycle.
  --             For each transfer between the FIFO register and the wr.axi_data_buffer, the counters of the number of bytes left of the 
  --             batch and the number of beats of the burst are decremented appropiatedly.
  -- Outside of 
  -- the FSM ->
  --         RD:A FIFO memory is used to store each beat transfered from the AXI read transaction, no matter from which subordinate.
  --            The BM transfer logic checks out if any more data is available from the RD FIFO to BM transfer, sending the data and 
  --            BM control signals bm_valid and bm_done. This last indicating the completion of the whole transaction at the last BM transfer.
  --            The BM transfer logic rearrenges the data to only transfer the data requested, even if the request is unaligned with 
  --            the AXI data bus width. This also includes applying a byte mask on the last BM transfer.
  --            Each BM transfer is done between the FIFO and the rd_burst.bm_data_buffer (which in between is the byte mask), so the BM 
  --            component connection has slack for a high fMAX synthesis. In addition, the rd_burst.bm_valid flag is high only when this 
  --            buffer contains valid data to be read by the BM component.
  --         WR:The wr.bm_data_buffer is used to read from the BM component the data to transfer in the write transaction.
  --            This is rearrenged and loaded into the FIFO register depending on the address it has been requested and how filled it is. 
  --            In case where the FIFO is full, the interface will deassert the wr.bm_ready so the bm_out.data_full is high.
  --            If there's not enough space on the present FIFO register, it will continue the write on the next. Due to this, it is 
  --            more efficient to have at least 4 registers on the WR FIFO, where on the RD FIFO it doesn't matter if it's 2 registers.
  --            
  --

  type rd_data_buffer   is array (natural range <>) of std_logic_vector( DATA_WIDTH - 1 downto 0 );
  type size_counter_arr is array (0 to 1) of unsigned(bm_in.rd_size'high + 1 downto 0);
  type main_state       is (idle, check_4kB, prepare_hs, handshake);
  type burst_state      is (idle, transfer, prepare_hs, handshake);

  -- Handshake type for read transactions. It's duplicated on rd_main and rd_burst to allow granting BM transactions while bursting.
  type rd_handshake_operation is record
    burst_4kb     : std_logic; -- Flag asserted when two bursts are required to complete the transaction due to surpassing the 4KB boundary.
    bm_size       : std_logic_vector(sel(12, 11, Mult_bursts_subor) downto 0);-- Original size being requested by BM component, and then first burst size.
    rem_size      : std_logic_vector(11 downto 0);-- Remaining size for second burst (4KB outbounds access)
    bm_addr       : std_logic_vector( ADDR_WIDTH     - 1 downto 0); -- Starting pointer requested by BM component.

    axi_mode      : std_logic_vector(1 downto 0); -- AXI output parameter: burst mode (FIXED, INC, WRAP).
    axi_cache     : std_logic_vector(3 downto 0); -- AXI output parameter: cache mode.
    axi_prot      : std_logic_vector(2 downto 0); -- AXI output parameter: privilage level access.
    axi_size      : std_logic_vector(2 downto 0); -- AXI output parameter: size mode of each beat in the burst.
    axi_len       : std_logic_vector(7 downto 0); -- AXI output parameter: number of beats in the burst.
    axi_addr      : std_logic_vector( ADDR_WIDTH     - 1 downto 0); -- AXI output parameter: Starting pointer of the AXI burst.
    axi_valid     : std_logic;                    -- AXI output parameter: valid flag for output control signals (addr, len, size, mode).

    start_shift   : unsigned( AXI4_DATA_BYTE - 1 downto 0); -- Number of right-bytes to skip when reading or writing data_bus at start of BM transfer.
    end_strb      : unsigned( AXI4_DATA_BYTE - 1 downto 0); -- Number of bytes to read from data_bus at the last BM transfer.
  end record rd_handshake_operation; 

  -- Initial handshake type for read transactions.
  type rd_main_operation is record
    state         : main_state;             -- State of the main handshake on read transactions.
    bm_grant      : std_logic;              -- Grant transaction request to BM component.
    hs            : rd_handshake_operation; -- Handshake control data to be AXI granted and sent to burst operation type.
  end record rd_main_operation;

  -- Burst type for read transactions.
  type rd_burst_operation is record
    state         : burst_state;            -- State of the read transaction.
    bm_error      : std_logic;              -- Error flag register due to SLVERR or DECERR subordinate response.

    hs            : rd_handshake_operation; -- Control data for AXI handshake
    axi_ready     : std_logic;              -- AXI output parameter: ready flag for input read data.

    fifo          : rd_data_buffer(   rd_n_fifo_regs - 1 downto 0); -- AXI data bus registers which filters narrow reads from data_tmp.
    fifo_full     : std_logic_vector( rd_n_fifo_regs - 1 downto 0); -- When asserted, the FIFO register is full or at a BM transfer.
    fifo_last     : std_logic_vector( rd_n_fifo_regs - 1 downto 0); -- When asserted, the FIFO register is the last BM transfer batch.

    bm_first      : std_logic;                                      -- Flag asserted until the first BM transfer has been done.
    bm_counter    : unsigned( AXI4_DATA_BYTE             downto 0); -- Used to count the number of bytes to BM transfer.
    bm_fifo_last  : std_logic;                                      -- BM transfers of the last AXI beat for the whole transaction flag.
    bm_valid      : std_logic;                                      -- Valid read data to transfer into BM bus from data_bus(dbits-1 downto 0).
    bm_done       : std_logic;                                      -- Asserted at the last rd_burst.bm_valid pulse of the whole transfer.

    bm_fifo_full      : std_logic_vector(rd_n_fifo_regs - 1 downto 0); -- fifo_full buffered register.
    data_fwidth       : std_logic_vector(DATA_WIDTH + dbits - 1 downto 0 ); -- Full shifted data bus
  end record rd_burst_operation;

  -- Handshake type for read transactions. It's duplicated on rd_main and rd_burst.
  type wr_handshake_operation is record
    burst_4kb     : std_logic; -- Flag asserted when two bursts are required to complete the transaction due to surpassing the 4KB boundary.
    bm_size       : std_logic_vector(sel(12, 11, Mult_bursts_subor) downto 0);-- Original size being requested by BM component, and then first burst size.
    rem_size      : std_logic_vector(11 downto 0);-- Remaining size for second burst (4KB outbounds access)
    bm_addr       : std_logic_vector( ADDR_WIDTH     - 1 downto 0); -- Starting pointer requested by BM component.

    axi_mode      : std_logic_vector(1 downto 0); -- AXI output parameter: burst mode (FIXED, INC, WRAP).
    axi_cache     : std_logic_vector(3 downto 0); -- AXI output parameter: cache mode.
    axi_prot      : std_logic_vector(2 downto 0); -- AXI output parameter: privilage level access.
    axi_size      : std_logic_vector(2 downto 0); -- AXI output parameter: size mode of each beat in the burst.
    axi_len       : std_logic_vector(7 downto 0); -- AXI output parameter: number of beats in the burst decremented by 1.
    axi_addr      : std_logic_vector( ADDR_WIDTH     - 1 downto 0); -- AXI output parameter: Starting pointer of the AXI burst.
    axi_strobe    : std_logic_vector( DATA_WIDTH/8   - 1 downto 0); -- AXI output parameter: What AXI data lanes to read from during AXI transfer.
    axi_valid     : std_logic;                    -- AXI output parameter: valid flag for output control signals (addr, len, size, mode).
  end record wr_handshake_operation; 

  type wr_main_operation is record
    state         : main_state;       -- State of the main handshake on write transactions.
    bm_grant      : std_logic;        -- Grant signals to BM component.
    hs            : wr_handshake_operation;
  end record wr_main_operation;

  type wr_burst_operation is record
    state         : burst_state;      -- State of the ongoing burst.
    bm_error      : std_logic;        -- Error flag register due to SLVERR or DECERR subordinate response.
    hs            : wr_handshake_operation;       -- Control data for AXI handshake.

    axi_valid_data: std_logic;                    -- AXI output parameter: valid write flag for output data.
    axi_first     : std_logic;                    -- First AXI beat of the burst flag used to compute the write strobe for that beat.

    fifo          : rd_data_buffer(   wr_n_fifo_regs - 1 downto 0); -- AXI data bus registers which filters narrow reads from data_tmp.
    fifo_full     : std_logic_vector( wr_n_fifo_regs - 1 downto 0); -- When asserted, the FIFO register is full or at a BM transfer.

    bm_active     : std_logic;                                      -- BM transfer active.
    bm_full_size  : unsigned(12 downto 0);                          -- BM size requested.
    bm_counter    : unsigned( AXI4_DATA_BYTE         - 1 downto 0); -- Used to count how many bytes have been filled on the actual FIFO register.

    bm_data_buffer : std_logic_vector( dbits         - 1 downto 0); -- BM data bus buffer, used to separate it from the BM component.
  end record wr_burst_operation;

  constant RST_RD_HANDSHAKE : rd_handshake_operation  := (
    burst_4kb         => '0',
    bm_size           => (others => '0'),
    rem_size          => (others => '0'),
    bm_addr           => (others => '0'),
    axi_mode          => "01",
    axi_cache         => (others => '0'),
    axi_prot          => (others => '0'),
    axi_size          => (others => '0'),
    axi_len           => (others => '0'),
    axi_addr          => (others => '0'),
    axi_valid         => '0',
    start_shift       => (others => '0'),
    end_strb          => (others => '0')
  );

  constant RST_RD_MAIN      : rd_main_operation       := (
    state             => idle,
    bm_grant          => '0',
    hs                => RST_RD_HANDSHAKE
  );

  constant RST_RD_BURST     : rd_burst_operation      := (
    state             => idle,
    bm_error          => '0',
    hs                => RST_RD_HANDSHAKE,
    axi_ready         => '0',
    fifo              => (others => (others => '0')),
    fifo_full         => (others => '0'),
    fifo_last         => (others => '0'),
    bm_first          => '1',
    bm_counter        => (others => '0'),
    bm_fifo_last      => '0',
    bm_valid          => '0',
    bm_done           => '0',
    bm_fifo_full      => (others => '0'),
    data_fwidth       => (others => '0')
  );

  constant RST_WR_HANDSHAKE : wr_handshake_operation  := (
    burst_4kb         => '0',
    bm_size           => (others => '0'),
    rem_size          => (others => '0'),
    bm_addr           => (others => '0'),
    axi_mode          => "01",
    axi_cache         => (others => '0'),
    axi_prot          => (others => '0'),
    axi_size          => (others => '0'),
    axi_len           => (others => '0'),
    axi_addr          => (others => '0'),
    axi_strobe        => (others => '0'),
    axi_valid         => '0'
  );

  constant RST_WR_MAIN      : wr_main_operation       := (
    state             => idle,
    bm_grant          => '0',
    hs                => RST_WR_HANDSHAKE
  );

  constant RST_WR_BURST     : wr_burst_operation      := (
    state             => idle,
    bm_error          => '0',
    hs                => RST_WR_HANDSHAKE,
    axi_valid_data    => '0',
    axi_first         => '1',
    fifo              => (others => (others => '0')),
    fifo_full         => (others => '0'),
    bm_active         => '0',
    bm_full_size      => (others => '0'),
    bm_counter        => (others => '0'),
    bm_data_buffer    => (others => '0')
  );

  -----------------------------------------------------------------------------
  -- Signal declaration
  -----------------------------------------------------------------------------

  -- Registers for write/read control.
  signal rd_main  : rd_main_operation;
  signal rd_burst : rd_burst_operation;
  signal wr_main  : wr_main_operation;
  signal wr_burst : wr_burst_operation;

  -- Handshake grant signals for main and burst loops for each transaction type.
  signal rd_main_axi_grant  : std_logic;
  signal rd_burst_axi_grant : std_logic;
  signal wr_burst_axi_grant : std_logic;
  signal wr_main_axi_grant  : std_logic;

  -- Injector mode registers.
  signal rd_size  : size_counter_arr;
  signal wr_size  : size_counter_arr;


  -----------------------------------------------------------------------------
  -- Function/procedure declaration
  -----------------------------------------------------------------------------

  -- To compute the number of beats required in the burst (length), the size requested is added to the LSB 
  -- of the starting address that has been requested. This sum contains the number of beats on the field 
  -- over AXI4_DATA_BYTE, since each beat use the whole AXI data bus width (DATA_WIDTH).
  function decide_len(
    bm_size   : std_logic_vector(MAX_BURST_BYTE - 1 downto 0);      -- Transfer size of the burst (real num needs +1)
    bm_addr   : std_logic_vector(rd_main.hs.bm_addr'high downto 0)  -- BM request address
  ) return std_logic_vector is 
      variable len_temp : std_logic_vector(MAX_BURST_BYTE - 1 downto 0);
  begin
    -- Number of bytes to AXI transfer (it cannot surpass 4kB) = BM address + BM size
    len_temp  := add_vector(bm_addr(AXI4_DATA_BYTE - 1 downto 0), bm_size, len_temp'length);

    -- If AXI DATA_WIDTH > 128 bits, the length will never surpass 256 (xFF), but requires padding with zeros.
    if(DATA_WIDTH > 128) then
      return (AXI4_DATA_BYTE + 7 downto MAX_BURST_BYTE => '0') & len_temp(MAX_BURST_BYTE - 1 downto AXI4_DATA_BYTE);
    -- If AXI DATA_WIDTH = 128 bits, the length will never surpass 256 (xFF), but it doesn't require padding.
    elsif(DATA_WIDTH = 128) then
      return len_temp(MAX_BURST_BYTE - 1 downto AXI4_DATA_BYTE);
    -- If AXI DATA_WIDTH < 128 bits, the length is on the MSB starting from AXI4_DATA_BYTE. However, if any bit 
    -- higher than AXI4_DATA_BYTE + 7 is asserted, the length will be 256 beats (xFF) and additional bursts will
    -- be necessary for this batch (thus, Mult_bursts_subor flag is TRUE).
    elsif(len_temp(MAX_BURST_BYTE downto AXI4_DATA_BYTE + 8) = (MAX_BURST_BYTE downto AXI4_DATA_BYTE + 8 => '0')) then
      return len_temp(AXI4_DATA_BYTE + 7 downto AXI4_DATA_BYTE);
    else
      return x"FF";
    end if;

  end function decide_len;

  
begin -- rtl

  -----------------
  -- Assignments --
  -----------------
  
  -- The assignments to the AXI interconnect bus are set in such way where the burst 
  -- handshake requests are prioritized over the ones requested by main.
  handshake_priority : process (rd_main, rd_burst, wr_main, wr_burst, axi4mi)
  begin
    -- Advance eXtensible Interface (interconnect bus)
      -- Write address channel out
    if(wr_burst.hs.axi_valid = '1') then
      axi4mo.aw_id      <= (axi4mo.aw_id'high   downto ID_W_WIDTH => '0') & std_logic_vector( to_unsigned(axi_id, ID_W_WIDTH) );
      axi4mo.aw_addr    <= (axi4mo.aw_addr'high downto ADDR_WIDTH => '0') & wr_burst.hs.axi_addr(ADDR_WIDTH-1 downto AXI4_DATA_BYTE) 
                          & (AXI4_DATA_BYTE-1 downto 0 => '0'); -- Address
      axi4mo.aw_region  <= (others => '0');
      axi4mo.aw_len     <= wr_burst.hs.axi_len;  -- Number of beats
      axi4mo.aw_size    <= wr_burst.hs.axi_size; -- Beat size
      axi4mo.aw_burst   <= wr_burst.hs.axi_mode; -- Burst mode
      axi4mo.aw_lock    <= '0';
      axi4mo.aw_cache   <= wr_burst.hs.axi_cache;
      axi4mo.aw_prot    <= wr_burst.hs.axi_prot;
      axi4mo.aw_qos     <= (others => '0');
      axi4mo.aw_valid   <= wr_burst.hs.axi_valid;
    elsif(rd_main.hs.axi_valid = '1') then -- TODO: DO AS SAME AS RD
      axi4mo.aw_id      <= (axi4mo.aw_id'high   downto ID_W_WIDTH => '0') & std_logic_vector( to_unsigned(axi_id, ID_W_WIDTH) );
      axi4mo.aw_addr    <= (axi4mo.aw_addr'high downto ADDR_WIDTH => '0') & wr_main.hs.axi_addr(ADDR_WIDTH-1 downto AXI4_DATA_BYTE) 
                          & (AXI4_DATA_BYTE-1 downto 0 => '0'); -- Address
      axi4mo.aw_region  <= (others => '0');
      axi4mo.aw_len     <= wr_main.hs.axi_len;  -- Number of beats
      axi4mo.aw_size    <= wr_main.hs.axi_size; -- Beat size
      axi4mo.aw_burst   <= wr_main.hs.axi_mode; -- Burst mode
      axi4mo.aw_lock    <= '0';
      axi4mo.aw_cache   <= wr_main.hs.axi_cache;
      axi4mo.aw_prot    <= wr_main.hs.axi_prot;
      axi4mo.aw_qos     <= (others => '0');
      axi4mo.aw_valid   <= wr_main.hs.axi_valid;
    else
      axi4mo.aw_id      <= (others => '0');
      axi4mo.aw_addr    <= (others => '0');
      axi4mo.aw_region  <= (others => '0');
      axi4mo.aw_len     <= (others => '0');
      axi4mo.aw_size    <= (others => '0');
      axi4mo.aw_burst   <= (others => '0');
      axi4mo.aw_lock    <= '0';
      axi4mo.aw_cache   <= (others => '0');
      axi4mo.aw_prot    <= (others => '0');
      axi4mo.aw_qos     <= (others => '0');
      axi4mo.aw_valid   <= '0';
    end if;
      -- Write data channel out
    axi4mo.w_data       <= (axi4mo.w_data'high downto DATA_WIDTH   => '0') & wr_burst.fifo(0);
    axi4mo.w_strb       <= (axi4mo.w_strb'high downto DATA_WIDTH/8 => '0') & wr_burst.hs.axi_strobe;
    --axi4mo.w_last       <= wr_burst.axi_last; -- Not registered, direct signalling
    axi4mo.w_valid      <= wr_burst.axi_valid_data;
      -- Write response channel out
    axi4mo.b_ready      <= '1';
      -- Read address channel out
    if(rd_burst.hs.axi_valid = '1') then
      axi4mo.ar_id      <= (axi4mo.ar_id'high   downto ID_R_WIDTH => '0') & std_logic_vector(to_unsigned(axi_id, ID_R_WIDTH));
      axi4mo.ar_addr    <= (axi4mo.ar_addr'high downto ADDR_WIDTH => '0') & rd_burst.hs.axi_addr(ADDR_WIDTH-1 downto AXI4_DATA_BYTE) 
                           & (AXI4_DATA_BYTE-1 downto 0 => '0'); -- Starting address
      axi4mo.ar_region  <= (others => '0');
      axi4mo.ar_len     <= rd_burst.hs.axi_len;  -- Number of beats
      axi4mo.ar_size    <= rd_burst.hs.axi_size; -- Beat size
      axi4mo.ar_burst   <= rd_burst.hs.axi_mode; -- Burst mode
      axi4mo.ar_lock    <= '0';
      axi4mo.ar_cache   <= rd_burst.hs.axi_cache;
      axi4mo.ar_prot    <= rd_burst.hs.axi_prot;
      axi4mo.ar_qos     <= (others => '0');
      axi4mo.ar_valid   <= rd_burst.hs.axi_valid;
    elsif(rd_main.hs.axi_valid = '1') then
      axi4mo.ar_id      <= (axi4mo.ar_id'high   downto ID_R_WIDTH => '0') & std_logic_vector(to_unsigned(axi_id, ID_R_WIDTH));
      axi4mo.ar_addr    <= (axi4mo.ar_addr'high downto ADDR_WIDTH => '0') & rd_main.hs.axi_addr(ADDR_WIDTH-1 downto AXI4_DATA_BYTE) 
                           & (AXI4_DATA_BYTE-1 downto 0 => '0'); -- Starting address
      axi4mo.ar_region  <= (others => '0');
      axi4mo.ar_len     <= rd_main.hs.axi_len;
      axi4mo.ar_size    <= rd_main.hs.axi_size;
      axi4mo.ar_burst   <= rd_main.hs.axi_mode;
      axi4mo.ar_lock    <= '0';
      axi4mo.ar_cache   <= rd_main.hs.axi_cache;
      axi4mo.ar_prot    <= rd_main.hs.axi_prot;
      axi4mo.ar_qos     <= (others => '0');
      axi4mo.ar_valid   <= rd_main.hs.axi_valid;
    else
      axi4mo.ar_id      <= (others => '0');
      axi4mo.ar_addr    <= (others => '0');
      axi4mo.ar_region  <= (others => '0');
      axi4mo.ar_len     <= (others => '0');
      axi4mo.ar_size    <= (others => '0');
      axi4mo.ar_burst   <= (others => '0');
      axi4mo.ar_lock    <= '0';
      axi4mo.ar_cache   <= (others => '0');
      axi4mo.ar_prot    <= (others => '0');
      axi4mo.ar_qos     <= (others => '0');
      axi4mo.ar_valid   <= '0';
    end if;
      -- Read data channel out
    axi4mo.r_ready      <= rd_burst.axi_ready;
      -- Write address channel in
    if(wr_burst.hs.axi_valid = '1') then
      wr_burst_axi_grant  <= axi4mi.aw_ready;
      wr_main_axi_grant   <= '0';
    elsif(wr_main.hs.axi_valid = '1') then
      wr_burst_axi_grant  <= '0';
      wr_main_axi_grant   <= axi4mi.aw_ready;
    else
      wr_burst_axi_grant  <= '0';
      wr_main_axi_grant   <= '0';
    end if;
      -- Write data channel in
    --axi4mi.w_ready; -- used as input
      -- Write response channel in
    --axi4mi.b_id;    -- used as input
    --axi4mi.b_resp;  -- used as input
    --axi4mi.b_valid; -- used as input
      -- Read address channel in
    if(rd_burst.hs.axi_valid = '1') then
      rd_burst_axi_grant  <= axi4mi.ar_ready;
      rd_main_axi_grant   <= '0';
    elsif(rd_main.hs.axi_valid = '1') then
      rd_burst_axi_grant  <= '0';
      rd_main_axi_grant   <= axi4mi.ar_ready;
    else
      rd_burst_axi_grant  <= '0';
      rd_main_axi_grant   <= '0';
    end if;
      -- Read data channel in
    --axi4mi.r_id;    -- used as input
    --axi4mi.r_data;  -- used as input
    --axi4mi.r_resp;  -- used as input
    --axi4mi.r_last;  -- used as input
    --axi4mi.r_valid; -- used as input

    -- Bus Master (injector)
      -- Write channel
    --bm_in.wr_addr;  -- used as input
    --bm_in.wr_size;  -- used as input
    --bm_in.wr_req;   -- used as input
    --bm_in.wr_data;  -- used as input
    bm_out.wr_req_grant <= wr_main.bm_grant;
    --bm_out.wr_full      <= not(wr_burst.bm_ready);  -- Not registered, direct signalling
    --bm_out.wr_done      <= wr_burst.bm_done;        -- Not registered, direct signalling
    bm_out.wr_err       <= wr_burst.bm_error;

      -- Read channel
    --bm_in.rd_addr;  -- used as input
    --bm_in.rd_size;  -- used as input
    --bm_in.rd_req;   -- used as input
    bm_out.rd_req_grant <= rd_main.bm_grant;
    bm_out.rd_data      <= (1023-dbits downto 0 => '0') & rd_burst.data_fwidth(dbits - 1 downto 0);
    bm_out.rd_valid     <= rd_burst.bm_valid;
    bm_out.rd_done      <= rd_burst.bm_done;
    bm_out.rd_err       <= rd_burst.bm_error;
  end process handshake_priority;
  
  -----------------------------------------------------------------------------
  -- Sequential process
  -----------------------------------------------------------------------------

  ------------------
  -- READ PROCESS --
  ------------------
  read_proc : process (clk, rstn) -- Variables used as connections between combinational logic, functions and registers.
    variable rd_addr_end          : std_logic_vector( 12             downto 0 );-- max end address LSB at INC mode (4kB check)

    variable rd_hs_done           : std_logic;                                  -- Flag to indicate the main handshake has been done.
    variable rd_burst_on          : std_logic;                                  -- Flag to start the burst transfer logic.
    variable rd_fifo_free_bottom  : std_logic;                                  -- Recursive flag to know if lower FIFO registers are free.
    variable rd_data_empty        : boolean;                                    -- rd.fifo(bm_index) register depleted flag. TODO: MAYBE ERASE THIS

    -- Variables only used on implementations where DATA_WIDTH < 128 bits.
    variable rd_next_bm_size      : std_logic_vector(rd_burst.hs.bm_size'range);-- Num of bytes left to transfer on the next clk cycle of this burst.

    -- Variables used only when injector mode is enabled. TODO: CLEAN THIS VAR IF NOT NECESSARY
    --variable size_threshold       : unsigned(AXI4_DATA_BYTE downto 0);
    
  begin
    if (rstn = '0' and ASYNC_RST) then
       -- Default variable values
      rd_main               <= RST_RD_MAIN;
      rd_burst              <= RST_RD_BURST;
      rd_hs_done            := '0';
      rd_burst_on           := '0';
      rd_fifo_free_bottom   := '0';
      rd_next_bm_size       := (others => '0');
      rd_size               <= (others => (others => '0'));
    elsif rising_edge(clk) then
      if (rstn = '0') then
        rd_main             <= RST_RD_MAIN;
        rd_burst            <= RST_RD_BURST;
        rd_hs_done          := '0';
        rd_burst_on         := '0';
        rd_fifo_free_bottom := '0';
        rd_next_bm_size     := (others => '0');
        rd_size             <= (others => (others => '0'));
      else
        -- Default var values
        rd_hs_done          := '0';
        rd_burst_on         := '0';
        rd_fifo_free_bottom := '0';
        rd_next_bm_size     := (others => '0');

        -- When injector mode is enabled, push new size if ongoing BM transfer finished.
        if(injector_mode and rd_size(0) = (rd_size'range => '0')) then
          rd_size(0) <= rd_size (1);
        end if;

        -----------------------------
        -- RD MAIN HANDSHAKE LOGIC --
        -----------------------------
        case rd_main.state is
          when idle =>
            -- Reset registers
            rd_main           <= RST_RD_MAIN;
            rd_main.bm_grant  <= '1';
          
            -- Load request information from BM
            if (bm_in.rd_req = '1' and rd_main.bm_grant = '1') then
              rd_main.bm_grant      <= '0'; -- Deassert granting requests for BM component
              rd_main.hs.bm_addr    <= bm_in.rd_addr(rd_main.hs.bm_addr'range); -- Load starting address request
              rd_main.hs.bm_size    <= (rd_main.hs.bm_size'high downto bm_in.rd_size'length => '0') & bm_in.rd_size; -- Size -1 from real
              rd_main.hs.axi_mode   <= '0' & not(bm_in.rd_fixed_addr);
              rd_main.hs.axi_cache  <= bm_in.rd_axi_cache;
              rd_main.hs.axi_prot   <= bm_in.rd_axi_prot;

              -- When injector mode is enabled, load real size on the queue.
              if(injector_mode) then
                rd_size(1)          <= unsigned('0' & bm_in.rd_size) + 1; -- Real size
              end if;

              -- Next, check 4kB out of bounds access
              rd_main.state         <= check_4kB;
            end if;
          
          
          when check_4kB =>
            -- Check if transaction will access two 4KB address regions
            rd_addr_end             := add_vector(rd_main.hs.bm_size, rd_main.hs.bm_addr(11 downto 0), rd_addr_end'length);
            rd_main.hs.burst_4kb    <= rd_addr_end(12);
          
            -- If transaction must be split in two bursts due to 4KB overflow boundary, calculate...
            if(rd_addr_end(12) = '1') then
              -- first burst size (-1 from real size)  MAX=4095, MIN=0
              rd_main.hs.bm_size    <= sub_vector(x"FFF", rd_main.hs.bm_addr(11 downto 0), rd_main.hs.bm_size'length);
              -- second burst size (-1 from real size) MAX=4094, MIN=0
              rd_main.hs.rem_size   <= rd_addr_end(rd_main.hs.rem_size'range);
            end if;
          
            -- Number of bytes to transfer at the last BM transfer = LSB ending address + 1 due to size being -1 from real
            rd_main.hs.end_strb     <= unsigned(rd_addr_end(AXI4_DATA_BYTE - 1 downto 0)) + 1;
          
            -- Next, compute size mode
            rd_main.state           <= prepare_hs;
          
          
          when prepare_hs =>
            -- Set AXI size mode to DATA_WIDTH and align the starting address with the DATA_WIDTH slot.
            rd_main.hs.axi_size     <= std_logic_vector(to_unsigned(AXI4_DATA_BYTE, rd_main.hs.axi_size'length));
            rd_main.hs.axi_addr     <= rd_main.hs.bm_addr(rd_main.hs.bm_addr'high downto AXI4_DATA_BYTE) & (AXI4_DATA_BYTE - 1 downto 0 => '0');

            -- Compute how many beats will be necessary to transfer the requested data in this burst.
            rd_main.hs.axi_len      <= decide_len(rd_main.hs.bm_size(11 downto 0), rd_main.hs.bm_addr);
          
            -- Save the number of bytes to discard unrequested data at the first BM transfer = LSB BM unaligned address + BM data bus width bytes
            rd_main.hs.start_shift  <= unsigned(rd_main.hs.bm_addr(AXI4_DATA_BYTE - 1 downto 0));
          
            -- Request AXI read burst when burst loop is on idle or bursting the last beat of the last burst. To verify the later when 
            -- Mult_bursts_subor = TRUE, an additional check must be performed (rd_burst.hs.bm_size < 256*DATA_WIDTH/8).
            if( rd_burst.state = idle 
            or(not(Mult_bursts_subor) and axi4mi.r_last = '1' and rd_burst.hs.burst_4kb = '0'           )
            or(    Mult_bursts_subor  and axi4mi.r_last = '1' and rd_burst.hs.burst_4kb = '0' 
                                      and rd_burst.hs.bm_size(rd_burst.hs.bm_size'high downto AXI4_DATA_BYTE + 8) 
                                          = (rd_burst.hs.bm_size'high downto AXI4_DATA_BYTE + 8 => '0') ) ) then
              rd_main.hs.axi_valid  <= '1';
              rd_main.state         <= handshake;
            end if;
            
          
          when handshake =>
            if( (rd_main_axi_grant and rd_main.hs.axi_valid) = '1') then
              rd_main.hs.axi_valid  <= '0'; -- At request being granted, deassert request
              rd_hs_done            := '1';
            end if;

            -- Once the burst is granted and the burst logic is on idle, send the control data to the burst logic.
            if(rd_burst.state = idle and (rd_main.hs.axi_valid = '0' or rd_hs_done = '1')) then
              rd_burst_on         := '1';
              rd_main             <= RST_RD_MAIN; -- Return idle to keep granting BM requests.
              rd_main.bm_grant    <= '1';
            end if;

        end case;
          
        -----------------------------
        -- RD BURST TRANSFER LOGIC --
        -----------------------------
        case rd_burst.state is
          when idle =>
            -- On command, initate the transfer of the burst.
            if(rd_burst_on = '1') then
              rd_burst.hs         <= rd_main.hs;-- Pass to burst the handshake control data.
              rd_burst.state      <= transfer;  -- Start transfering data
              rd_burst.axi_ready  <= '1';
            end if;

          when transfer => -- AXI transfer --
          -- The AXI transfer occurs by buffering the read data onto the rd_burst.axi_data_buffer register when the subordinate asserts the valid data flag.
          -- Then, the rd_burst.axi_data_buffer is loaded onto a FIFO register, which will be used at the BM transfer. However, due to this single clock 
          -- cycle delay between AXI read and data load, both valid and the mask signals are also buffered on the "buffer" registers (these
          -- are outside of the state machine and updated with each clock pulse). 

              -- Check if subordinate is delivering valid data with the same AXI ID as requested and if manager is listening.
            if (axi4mi.r_valid = '1' and axi4mi.r_id(ID_R_WIDTH-1 downto 0) = std_logic_vector(to_unsigned(axi_id, ID_R_WIDTH)) 
                and rd_burst.axi_ready = '1') then

              -- Register inputs to separate AXI network from further computation.
              rd_burst.fifo(rd_n_fifo_regs - 1) <= axi4mi.r_data(DATA_WIDTH - 1 downto 0);
              rd_burst.bm_error                 <= axi4mi.r_resp(1);

              -- Signal the present rd_burst.FIFO register as prepared for BM transfer, for whenever it is due to FIFO queue.
              rd_burst.fifo_full(rd_n_fifo_regs - 1)   <= '1';

              -- Deassert the ready flag to finish the AXI burst if it is the last beat or if there is not enough space in the FIFO at the moment.
              if( axi4mi.r_last = '1' or rd_burst.fifo_full(rd_n_fifo_regs - 2 downto 0) = (rd_n_fifo_regs - 2 downto 0 => '1') ) then
                rd_burst.axi_ready    <= '0';
              end if;

              -- The last AXI transfer of the whole transaction will set the proper rd_burst.fifo_last bit, so the BM transfer logic knows when to end.
              -- However, there's a distinction between DATA_WIDTH <= 64 bits and higher data widths. If there's still data to transfer to the same 
              -- subordinate because this burst has not been enough, do not assert the last BM transfer on the FIFO register and update rd_burst.bm_size.
              if(Mult_bursts_subor) then
                rd_next_bm_size     := sub_vector(rd_burst.hs.bm_size, DATA_WIDTH/8, rd_next_bm_size'length);
                rd_burst.hs.bm_size <= rd_next_bm_size;
                -- Mark as last FIFO register to be read by BM if there is not another burst due to 4kB surpass, the last beat has been
                -- received as last of the burst and there's no more data for this burst (rd_next_bm_size is overflown due to the subtraction).
                rd_burst.fifo_last(rd_n_fifo_regs - 1)  <= not(rd_burst.hs.burst_4kb) and axi4mi.r_last and rd_next_bm_size(rd_next_bm_size'high);
              else
                rd_burst.fifo_last(rd_n_fifo_regs - 1)  <= not(rd_burst.hs.burst_4kb) and axi4mi.r_last;
              end if;

              -- On last AXI beat...
              if(axi4mi.r_last = '1') then
                -- Compute new handshake if multiple bursts are necessary to complete this data batch:
                if( Mult_bursts_subor and rd_next_bm_size(rd_next_bm_size'high) = '0' ) then
                  if(rd_burst.hs.axi_mode = INC) then
                    rd_burst.hs.axi_addr  <= add_vector(rd_burst.hs.axi_addr(rd_burst.hs.bm_addr'high downto 8 + AXI4_DATA_BYTE), 1, 
                                            rd_burst.hs.axi_addr'high - 7 - AXI4_DATA_BYTE) & (7 + AXI4_DATA_BYTE downto 0 => '0');
                  end if;
                  rd_burst.state          <= prepare_hs;

                -- Or compute a new handshake if there's another batch of data due to the 4kB split. 
                elsif(rd_burst.hs.burst_4kb = '1') then
                  if(Mult_bursts_subor) then
                    rd_burst.hs.bm_size   <= '0' & rd_burst.hs.rem_size;
                  else
                    rd_burst.hs.bm_size   <= rd_burst.hs.rem_size;
                  end if;
                  if(rd_burst.hs.axi_mode = INC) then
                    rd_burst.hs.axi_addr  <= add_vector(rd_burst.hs.axi_addr(rd_burst.hs.axi_addr'high downto 12), 1, 
                                               rd_burst.hs.axi_addr'high - 11) & (11 downto 0 => '0');
                  end if;
                  rd_burst.state          <= prepare_hs;
                else
                -- The transaction has finished on the AXI side.
                  rd_burst.state      <= idle;
                end if;
              end if;
            -- In case no read is happening, assert AXI ready if there's free space on the FIFO.
            elsif( (rd_burst.fifo_full(rd_n_fifo_regs - 2 downto 0) /= (rd_n_fifo_regs - 2 downto 0 => '1')) ) then
              rd_burst.axi_ready      <= '1';
            end if;


          when prepare_hs =>
            -- Compute how many beats will be necessary to transfer the requested data in this burst.
            rd_burst.hs.axi_len       <= decide_len(rd_burst.hs.bm_size(11 downto 0), rd_burst.hs.axi_addr);
          
            -- Next, the handshake step.
            rd_burst.hs.axi_valid     <= '1'; -- Request AXI read burst.
            rd_burst.state            <= handshake;


          when handshake =>
            -- Request burst transaction with priority over main loop.
            if( (rd_burst_axi_grant and rd_burst.hs.axi_valid) = '1') then
              rd_burst.hs.axi_valid   <= '0'; -- At request being granted, deassert request.
              -- Clean the 4kB flag when all burst of the same subordinate have finished.
              if( not(Mult_bursts_subor and rd_burst.hs.bm_size(rd_burst.hs.bm_size'high) /= '1') ) then
                rd_burst.hs.burst_4kb <= '0';
              end if;
              rd_burst.state          <= transfer;
            end if;

        end case;


      -------------------------
      -- RD BM DATA TRANSFER --
      -------------------------
        -- WIP: Due to technical difficulties that must be solved in the future, the BM transfer logic must be revised.
        --      Thus, for the moment, use the injector_mode that simulates the correct number of readings.
      -- The injector mode, when enabled, discards all read data while simulates the correct BM signaling for the transaction.
        if(injector_mode) then
          rd_burst.fifo_full(0) <= '0';
          rd_burst.fifo_last(0) <= '0';
          rd_fifo_free_bottom   := '1';
          rd_burst.bm_valid     <= '0';
          rd_burst.bm_done      <= '0';
          if(rd_size(0) /= (rd_size(0)'range => '0')) then
            rd_burst.bm_valid   <= '1';
            rd_size(0)          <= rd_size(0) - dbits/8;
            if(rd_size(0) <= dbits/8) then
              rd_burst.bm_done  <= '1';
              rd_size(0)        <= (others => '0');
            end if;
          end if;

        else -- INJECTOR_MODE = FALSE

      -- The BM transfer logic transfers from the RD FIFO to the BM component at dbits bits per clock cycle throughput without pause, unless  
      -- there's not enough data in the FIFO to BM transfer. This is achieved by loading rd_burst.fifo(bm_index) onto rd_burst.data_fwidth 
      -- used as output, which transfers data and shifts while there's enough to perform a BM transfer (rd_burst.bm_counter >= dbits/8). 
      -- When the rd_burst.data_fwidth does not have enough data for a BM transfer, the next FIFO register is read and positioned after the  
      -- data left to be read, freeing the FIFO register since it has been read for new AXI beat readings.

--          -- Set combinational variables --
--          -- Check if this is the last BM transfer before rd_burst.fifo(bm_index) is depleted after a transfer of dbits bits.
--          rd_data_empty       := rd_burst.bm_counter < to_unsigned(dbits/8, rd_burst.bm_counter'length);
--
--          -- Check if there's data to BM transfer. Delayed with a buffer register so the last AXI beat transfer is finished on this FIFO register.
--          if(rd_burst.bm_fifo_full(0) = '1' or rd_burst.bm_first = '0') then
--
--          -- Before any BM transfer, load and shift the FIFO register to put the requested data on 0 to higher, flushing unrequested data read 
--          -- by the AXI side. Then, initilize the rd_burst.bm_counter with [the whole AXI data bus width bytes value or with the number of bytes
--          -- to read from the last FIFO register to BM transfer] minus the shift performed on this rd_burst.bm_first cycle.
--            if(rd_burst.bm_first = '1') then
--
--              -- Deassert the first BM transfer flag, since it's only required to shift rd_burst.start_shift before than the first BM transfer.
--              rd_burst.bm_first   <= '0';
--
--              -- The initial counter is set by rd_burst.end_strb if there's only one FIFO register to transfer. 
--              if(rd_burst.fifo_last(0) = '1') then
--                rd_burst.bm_counter <= rd_burst.hs.end_strb - rd_burst.hs.start_shift;
--              else -- Otherwise, the initial counter is the AXI data bus bytes.
--                rd_burst.bm_counter <= to_unsigned(DATA_WIDTH/8, rd_burst.bm_counter'length) - rd_burst.hs.start_shift;
--              end if;
--
--              -- Load, shift and free the FIFO register. Also, record if this is the last AXI beat of the whole BM transaction.
--              rd_burst.data_fwidth  <= (rd_burst.data_fwidth'high downto DATA_WIDTH - 8*to_integer(rd_burst.hs.start_shift) => '0') 
--                                       & rd_burst.fifo(0)(DATA_WIDTH - 1 downto DATA_WIDTH - 8*to_integer(rd_burst.hs.start_shift));
--              rd_burst.fifo_full(0) <= '0';
--              rd_fifo_free_bottom   := '1';
--              rd_burst.bm_fifo_last <= rd_burst.fifo_last(0);
--
--          else -- rd_burst.bm_first = '0' check
--            if(not rd_data_empty) then
--
--              -- There's enough data to BM transfer on the next cycle, so shift a BM transfer.
--              rd_burst.data_fwidth  <= std_logic_vector(shift_right(unsigned(rd_burst.data_fwidth), dbits/8));
--
--              -- Update BM counter.
--              rd_burst.bm_counter   <= rd_burst.bm_counter - dbits/8;
--
--            else  -- There isn't enough data on rd_burst.data_fwidth to BM transfer.
--
--              -- Last BM transfer
--              if(rd_burst.bm_fifo_last = '1') then
--                -- TODO: Apply a mask, both in here and on the first BM transfer.
--                rd_burst.data_fwidth  <= (rd_burst.data_fwidth'high downto dbits => '0') & rd_burst.data_fwidth(dbits - 1 downto 0);
--                rd_burst.bm_counter   <= (others => '0');
--                rd_burst.bm_first     <= '1';
--
--              elsif(rd_burst.bm_fifo_full(0) = '1' or rd_burst.bm_fifo_last = '1') then
--
--              -- In case this cycle will deplete rd_burst.data_fwidth and the next FIFO register is prepared to be transfered,
--              -- use the remaining data (rd_burst.bm_counter lower or equal to AXI data bus bytes) as LSB and take the 
--              -- lacking bytes to fill dbits from the next FIFO register, while also shifting its content for posterior transfers.
--              -- (since the shifting index k surpasses the bytes available in the next FIFO register on unaligned starting transfers, 
--              -- fill the remaining byte positions with zeros, that, in number of bytes, will be always lower than the bytes in dbits)
--                rd_burst.data_fwidth  <= (DATA_WIDTH + 8*to_integer(rd_burst.bm_counter) - 1 downto dbits => '0') 
--                                          & rd_burst.fifo(0) 
--                                          & rd_burst.data_fwidth(8*to_integer(rd_burst.bm_counter) - 1 downto dbits);
--
--                -- Set the present FIFO register to be prepared for new AXI transfer and change the FIFO register rd_burst.bm_index.
--                rd_burst.fifo_full(0) <= '0';
--
--                -- Compute the number of bytes that'll be left to read on the next FIFO register.
--                -- In case where the next FIFO register is the last, counter = end_strb - ( dbits/8 - bm_counter ) = ( end_strb + bm_counter ) - dbits/8
--                -- Otherwise, it must be taken the whole AXI data bus, counter = AXI_DATA/8 - ( dbits/8 - bm_counter ) = bm_counter + AXI_DATA/8 - dbits/8
--                if(rd_burst.fifo_last(1) = '1') then
--                  rd_burst.bm_counter <= rd_burst.hs.end_strb + rd_burst.bm_counter - dbits/8;
--
--                  -- In addition, if the number of bytes read on this clock cycle from rd_burst.fifo(rd_bm_next_index) include all the data required 
--                  -- by rd_burst.end_strb, end the transfer on the next clock cycle. (done, mask and return to idle)
--                  if(to_unsigned(dbits/8, rd_burst.bm_counter'length) - rd_burst.bm_counter >= rd_burst.hs.end_strb) then
--                    rd_burst.bm_done  <= '1';
--                    rd_burst.state    <= idle;
--                  end if;
--
--                else
--                  rd_burst.bm_counter <= rd_burst.bm_counter + DATA_WIDTH/8 - dbits/8;
--                end if;              
--
--              else   -- rd_burst.fifo_full(rd_bm_next_index) = 0 check
--
--              -- In case there's not enough data to read from the FIFO, check if this is the last FIFO register to BM transfer. If it 
--              -- is, check how many bytes of remaining data are left. If it's lower than dbits/8, this is the last BM transfer. However, 
--              -- if it's exactly dbits/8 and it's the last FIFO register, delay the end of the BM transfer for another clock cycle 
--              -- (do not increase the rd_burst.bm_counter, let the execution return to this step to execute the end of the BM transfer).
--                if(rd_burst.fifo_last(0) = '1') then 
--                  rd_burst.bm_counter <= rd_burst.bm_counter - dbits/8;
--                  rd_burst.bm_done  <= '1';
--                  rd_burst.state    <= idle;
--                else
--              -- Otherwise, if there's not enough data and this is not the last FIFO register, wait for the next AXI transfer.
--                end if;
--
--              end if; -- rd_burst.fifo_full(rd_bm_next_index) end of check
--            end if; -- rd_empty_data end of check
--          end if;   -- bm_first end of check
--
--          if(rd_burst.bm_counter >= 2*dbits/8 or rd_burst.bm_fifo_last = '1' or rd_burst.bm_fifo_full(0) = '1' ) then
--            rd_burst.bm_valid     <= '1';
--          else
--            rd_burst.bm_valid     <= '0';
--          end if;
--
        end if; -- INJECTOR_MODE CHECK


        -- Delayed signals, to be revised.
        rd_burst.bm_fifo_full <= rd_burst.fifo_full;
        

      -------------
      -- RD FIFO --
      -------------
        -- On each clock cycle, push new data from top to the bottom on the FIFO, if bottom is or will be free.
        for k in 1 to rd_n_fifo_regs - 1 loop
          rd_fifo_free_bottom := rd_burst.fifo_full(k - 1) or rd_fifo_free_bottom;
          if(rd_fifo_free_bottom = '0') then
            rd_burst.fifo_full(k)     <= '0';
            rd_burst.fifo_full(k - 1) <= rd_burst.fifo_full(k);
            rd_burst.fifo_last(k - 1) <= rd_burst.fifo_last(k);
            rd_burst.fifo(k - 1)      <= rd_burst.fifo(k);
          end if;
        end loop;

      end if;
    end if;
  end process read_proc;



  -------------------
  -- WRITE PROCESS --
  -------------------
  write_proc : process (clk, rstn) -- Variables used as connections between combinational logic, functions and registers.
    variable wr_bm_start          : std_logic;                                      -- Start BM transfer
    variable wr_addr_end          : std_logic_vector( 12               downto 0 );  -- max end address LSB at INC mode (4kB check)
    variable wr_hs_done           : std_logic;                                      -- Flag to indicate the main handshake has been done.
    variable wr_fifo_free_bottom  : std_logic;                                      -- Free of the FIFO bottom

    -- Variables only used on implementations where DATA_WIDTH < 128 bits.
    variable wr_next_bm_size      : std_logic_vector(wr_burst.hs.bm_size'range);-- Num of bytes left to transfer on the next clk cycle of this burst.
    
  begin
    if (rstn = '0' and ASYNC_RST) then
      wr_main               <= RST_WR_MAIN;
      wr_burst              <= RST_WR_BURST;
      wr_bm_start           := '0';
      wr_addr_end           := (others => '0');
      wr_hs_done            := '0';
      wr_fifo_free_bottom   := '0';
    elsif rising_edge(clk) then
      if (rstn = '0') then
        wr_main             <= RST_WR_MAIN;
        wr_burst            <= RST_WR_BURST;
        wr_bm_start         := '0';
        wr_addr_end         := (others => '0');
        wr_hs_done          := '0';
        wr_fifo_free_bottom := '0';
      else
        wr_bm_start         := '0';
        wr_addr_end         := (others => '0');
        wr_hs_done          := '0';
        wr_fifo_free_bottom := '0';

      -----------------------------
      -- WR MAIN HANDSHAKE LOGIC --
      -----------------------------
        case wr_main.state is
          when idle =>
            -- Grant BM if previous BM transaction has been completed.
            wr_main.bm_grant        <= not(wr_burst.bm_active);
          
            -- Load request information from BM
            if (bm_in.wr_req = '1' and wr_main.bm_grant = '1') then
              wr_main.bm_grant      <= '0';           -- Deassert granting requests for BM component
              wr_main.hs.bm_addr    <= bm_in.wr_addr(wr_main.hs.bm_addr'range); -- Load starting address request
              wr_main.hs.bm_size    <= (wr_main.hs.bm_size'high downto bm_in.wr_size'length => '0') & bm_in.wr_size; -- Size -1 from real
              wr_main.hs.axi_mode   <= '0' & not(bm_in.wr_fixed_addr);
              wr_main.hs.axi_cache  <= bm_in.wr_axi_cache;
              wr_main.hs.axi_prot   <= bm_in.wr_axi_prot;

              -- Start the BM transfer on the next clock cycle.
              wr_burst.bm_active    <= '1';
              wr_bm_start           := '1';
              wr_burst.bm_full_size <= ((wr_burst.bm_full_size'high downto bm_in.wr_size'length => '0') & unsigned(bm_in.wr_size)) + 1; -- Real size

              -- Next, check 4kB out of bounds access
              wr_main.state         <= check_4kB;
            end if;
          
          
          when check_4kB => -- Worst delay path: ADD 12+12, SUB 13-13
            -- Check if transaction will access two 4KB address regions
            wr_addr_end             := add_vector(wr_main.hs.bm_size, wr_main.hs.bm_addr(11 downto 0), wr_addr_end'length);
            wr_main.hs.burst_4kb    <= wr_addr_end(12);
          
            -- If transaction must be split in two bursts, due to 4KB overflow boundary, calculate...
            if(wr_addr_end(12) = '1') then
              -- first burst size  (-1 from real size) MAX=4095, MIN=0
              wr_main.hs.bm_size    <= sub_vector(x"FFF", wr_main.hs.bm_addr(11 downto 0), wr_main.hs.bm_size'length);
              -- second burst size (-1 from real size) MAX=4094, MIN=0
              wr_main.hs.rem_size   <= wr_addr_end(wr_main.hs.rem_size'range);
            end if;

            -- Next, compute size mode
            wr_main.state           <= prepare_hs;
          
          
          when prepare_hs =>
            -- Set AXI size mode to DATA_WIDTH and align the starting address with the DATA_WIDTH slot.
            wr_main.hs.axi_size     <= std_logic_vector(to_unsigned(AXI4_DATA_BYTE, wr_main.hs.axi_size'length));
            wr_main.hs.axi_addr     <= wr_main.hs.bm_addr(wr_main.hs.bm_addr'high downto AXI4_DATA_BYTE) & (AXI4_DATA_BYTE - 1 downto 0 => '0');

            -- Compute how many beats will be necessary to transfer the requested data in this burst.
            wr_main.hs.axi_len      <= decide_len(wr_main.hs.bm_size(11 downto 0), wr_main.hs.bm_addr);

            -- Generate the mask to be shifted for the first AXI transfer.
            for k in wr_main.hs.axi_strobe'range loop
              if(k > to_integer(unsigned(wr_main.hs.bm_size(AXI4_DATA_BYTE - 1 downto 0)))) then
                wr_main.hs.axi_strobe(k) <= '0';
              else
                wr_main.hs.axi_strobe(k) <= '1';
              end if;
            end loop;
            
            -- Request AXI write burst when burst loop is on idle or bursting the last beat of the last burst. To verify the later when 
            -- Mult_bursts_subor = TRUE, an additional check must be performed (wr_burst.hs.bm_size < DATA_WIDTH).
            if( wr_burst.state = idle 
            or(not(Mult_bursts_subor) and wr_burst.hs.burst_4kb = '0'                                   ) 
            or(    Mult_bursts_subor  and wr_burst.hs.burst_4kb = '0' 
                                      and wr_burst.hs.bm_size(wr_burst.hs.bm_size'high downto AXI4_DATA_BYTE + 8) 
                                          = (wr_burst.hs.bm_size'high downto AXI4_DATA_BYTE + 8 => '0') ) ) then
              wr_main.hs.axi_valid      <= '1'; -- Request AXI write burst.
              wr_main.state             <= handshake;
            end if;
          
          
          when handshake =>
            -- Having all computation steps and proper registration separated allows maximum 
            -- frequency of operation when including this AXI manager interface at the interconnect
            -- bus. For a write burst, AW AXI control buses are used to send the burst control data.
            if (wr_main_axi_grant = '1' and wr_main.hs.axi_valid = '1') then
              wr_main.hs.axi_valid      <= '0'; -- At request being granted, deassert AXI handshake request.
              wr_hs_done                := '1';
            end if;

            if(wr_burst.state = idle and (wr_main.hs.axi_valid = '0' or wr_hs_done = '1')) then
              wr_burst.hs               <= wr_main.hs;
              -- Shift the initial mask and load it on the burst logic.
              wr_burst.hs.axi_strobe    <= std_logic_vector(shift_left( unsigned((wr_burst.hs.axi_strobe)), 
                                           to_integer(unsigned(wr_main.hs.bm_addr(AXI4_DATA_BYTE - 1 downto 0))) ));
              -- Add bm_address to first batch size so it's aligned with DATA_WIDTH. This, will be used as last beat strobe.
              wr_burst.hs.bm_size       <= add_vector(wr_main.hs.bm_size, wr_main.hs.bm_addr(AXI4_DATA_BYTE - 1 downto 0), 
                                           wr_burst.hs.bm_size'length);
              wr_burst.state            <= transfer;
              if(injector_mode) then
                wr_burst.axi_valid_data <= '1';
              else
                wr_burst.axi_valid_data <= wr_burst.fifo_full(1) or wr_burst.fifo_full(0);
              end if;
              
              -- Next, beat transfers
              wr_main.state             <= idle;
            end if;

        end case;


      -----------------------------
      -- WR BURST TRANSFER LOGIC --
      -----------------------------
        case wr_burst.state is 
          when idle =>
            null;


          when transfer => -- AXI transfer --
          -- The AXI transfer sets the AXI valid write flag anytime there's data available in a buffer register that reads from the FIFO, 
          -- freeing the FIFO register for BM fransfers. In addition, the size left to transfer wr.bm_size is decreased with the number of 
          -- bytes transfered.

            -- Load the variables for last AXI beat in the burst, next FIFO index at the AXI side and the read flag.
            wr_fifo_free_bottom           := wr_burst.axi_valid_data and axi4mi.w_ready;
            wr_burst.fifo_full(0)         <= wr_fifo_free_bottom;

            -- On the first beat read, zero the wr.bm_addr LSB used to set up the lower bound of the strobe for the first beat.
            -- Generate the mask to be shifted for the first AXI transfer.
            for k in wr_burst.hs.axi_strobe'range loop
              if(k > to_integer(unsigned(wr_burst.hs.bm_size(AXI4_DATA_BYTE - 1 downto 0)))) then
                wr_burst.hs.axi_strobe(k) <= '0';
              else
                wr_burst.hs.axi_strobe(k) <= '1';
              end if;
            end loop;

            -- Each AXI transfer, update size left on this batch.
            if(wr_fifo_free_bottom = '1') then
              wr_next_bm_size             := sub_vector(wr_burst.hs.bm_size, DATA_WIDTH/8, wr_burst.hs.bm_size'length);
              wr_burst.hs.bm_size         <= wr_next_bm_size;
              if(not(injector_mode)) then
                wr_burst.axi_valid_data   <= wr_burst.fifo_full(1);
              end if;

              -- Check if it's the last beat.
              if(wr_burst.hs.axi_len = (wr_burst.hs.axi_len'range => '0')) then
                axi4mo.w_last             <= '1';
                -- If multiple bursts to same subordinate may be necessary, check for those cases.
                if(Mult_bursts_subor and wr_next_bm_size(wr_next_bm_size'high) = '0') then
                    if(wr_burst.hs.axi_mode = INC) then
                      wr_burst.hs.axi_addr <= add_vector(wr_burst.hs.axi_addr(wr_burst.hs.bm_addr'high downto 8 + AXI4_DATA_BYTE), 1, 
                                                 wr_burst.hs.axi_addr'high - 7 - AXI4_DATA_BYTE) & (7 + AXI4_DATA_BYTE downto 0 => '0');
                    end if;
                    wr_burst.state        <= prepare_hs;
                -- If second burst/batch must be processed.
                elsif(wr_burst.hs.burst_4kb = '1') then
                  if(Mult_bursts_subor) then
                    wr_burst.hs.bm_size   <= '0' & wr_burst.hs.rem_size;
                  else
                    wr_burst.hs.bm_size   <= wr_burst.hs.rem_size;
                  end if;
                  if(wr_burst.hs.axi_mode = INC) then
                    wr_burst.hs.axi_addr  <= add_vector(wr_burst.hs.axi_addr(wr_burst.hs.axi_addr'high downto 12), 1, 
                                             wr_burst.hs.axi_addr'high - 11) & (11 downto 0 => '0');
                  end if;
                  wr_burst.state          <= prepare_hs;
                else
                -- Whole transaction has finished, return to idle.
                  wr_burst.state          <= idle;
                end if;
              end if;
            elsif(not(injector_mode)) then 
            -- No AXI beat has occured, check if there's data on the FIFO.
              wr_burst.axi_valid_data     <= wr_burst.fifo_full(0);
            end if;


          when prepare_hs =>
            -- Compute how many beats will be necessary to transfer the requested data in this burst.
            wr_burst.hs.axi_len           <= decide_len(wr_burst.hs.bm_size(11 downto 0), wr_burst.hs.axi_addr);
            wr_burst.hs.axi_valid         <= '1'; -- Request AXI write burst.

            wr_burst.state                <= handshake;


          when handshake =>
            -- Request burst transaction with priority over main loop.
            if( (wr_burst_axi_grant and wr_burst.hs.axi_valid) = '1') then
              wr_burst.hs.axi_valid       <= '0'; -- At request being granted, deassert request.
              -- Clean the 4kB flag when all burst of the same subordinate have finished.
              if( not(Mult_bursts_subor and wr_burst.hs.bm_size(wr_burst.hs.bm_size'high) /= '1') ) then
                wr_burst.hs.burst_4kb     <= '0';
              end if;
              if(injector_mode) then
                wr_burst.axi_valid_data   <= '1';
              else
                wr_burst.axi_valid_data   <= wr_burst.fifo_full(1) or wr_burst.fifo_full(0);
              end if;
              wr_burst.state              <= transfer;
            end if;


        end case;


      -------------------------
      -- WR BM DATA TRANSFER --
      -------------------------
        if(injector_mode) then
          if(wr_burst.bm_active = '1' or wr_bm_start = '1') then
            bm_out.wr_full              <= wr_burst.fifo_full(wr_n_fifo_regs - 2) and not(wr_fifo_free_bottom);
            if(wr_burst.bm_full_size > dbits/8) then
              wr_burst.bm_full_size     <= wr_burst.bm_full_size - dbits/8;
            else
              wr_burst.bm_full_size     <= (others => '0');
              bm_out.wr_done            <= '1';
              wr_burst.bm_active        <= '0';
            end if;
          else
            bm_out.wr_done              <= '0';
            bm_out.wr_full              <= '1';
          end if;
        else
          -- TODO: BUFFER BM DATA INPUT, REARRANGE AND PUT IT ON THE FIFO'S TOP
        end if;


      -------------
      -- WR FIFO --
      -------------
        -- On each clock cycle, push new data from top to the bottom on the FIFO, if bottom is or will be free.
        for k in 1 to wr_n_fifo_regs - 1 loop
          wr_fifo_free_bottom := wr_burst.fifo_full(k - 1) or wr_fifo_free_bottom;
          if(wr_fifo_free_bottom = '0') then
            wr_burst.fifo_full(k)     <= '0';
            wr_burst.fifo_full(k - 1) <= wr_burst.fifo_full(k);
            wr_burst.fifo(k - 1)      <= wr_burst.fifo(k);
          end if;
        end loop;

      -------------------------
      -- WRITE RESPONSE READ --
      -------------------------

        -- This logic always listen for write responses, not matter if a write transaction is not ongoing.
        if(axi4mi.b_valid = '1' and axi4mi.b_id(ID_W_WIDTH-1 downto 0) = std_logic_vector(to_unsigned(axi_id, ID_W_WIDTH))) then
          wr_burst.bm_error <= axi4mi.b_resp(1);
        end if;
      
      
      end if;
    end if;
  end process write_proc;

  -----------------------------------------------------------------------------
  -- Combinational process
  -----------------------------------------------------------------------------


end architecture rtl;